------------------------------------------------------------------------------
-- Strucutral description of a pipeline stage
------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE work.dxp_package.all;
------------------------------------------------------------------------------
entity dxp_PSLM_stage_vhdl is
	port (mr_Din					:	in		std_logic_vector(3 downto 0);
			Md_Din, FP_Din			:	in		std_logic_vector(7 downto 0);
			Clock, Reset, LD_All	:	in 	std_logic;
			mr_shr_out				:	out	std_logic_vector(3 downto 0);
			Md_shl_out, PP_out	:	out 	std_logic_vector(7 downto 0));
end dxp_PSLM_stage_vhdl;

architecture structural of dxp_PSLM_stage_vhdl is	
------------------------------------------------------------------------------			
signal and_out, Md_Dout, FP_Dout : std_logic_vector(7 downto 0);
signal mr_Dout : std_logic_vector(3 downto 0);
signal mrSDoutR, mrSDoutL, MdSDoutR, MdSDoutL, FPSDoutR, FPSDoutL : std_logic;
begin
------------------------------------------------------------------------------
-- The registers
------------------------------------------------------------------------------
mr_Reg :	dxp_nBitSFR_vhdl 	generic map (n => 4) 
	port map (mr_Din, '0', '0', Clock, Reset, LD_All, '0', '0', 
									mrSDoutR, mrSDoutL, mr_Dout);
Md_Reg :	dxp_nBitSFR_vhdl 	generic map (n => 8) 
	port map (Md_Din, '0', '0', Clock, Reset, LD_All, '0', '0', 
									MdSDoutR, MdSDoutL, Md_Dout);
FP_Reg :	dxp_nBitSFR_vhdl	generic map (n => 8) 
	port map (FP_Din, '0', '0', Clock, Reset, LD_All, '0', '0', 
									FPSDoutR, FPSDoutL, FP_Dout);
-------------------------------------------------------------------------------
-- Instead of the MUX in the SSLM, I use here a BIT-WISE AND. The left operand 
-- is generated by using the replication operator, i.e. it replicates 
-- mr_Dout[0] 8 times.
-------------------------------------------------------------------------------
	and_out <= (mr_Dout(0) & mr_Dout(0) & mr_Dout(0) & mr_Dout(0) & 
				mr_Dout(0) & mr_Dout(0) & mr_Dout(0) & mr_Dout(0)) and Md_Dout;
-------------------------------------------------------------------------------
-- The stage output assignments
-------------------------------------------------------------------------------
	PP_out <= and_out + FP_Dout; --You have to instantiate your adder here!!!
	mr_shr_out <= ('0' & mr_Dout(3 downto 1));
	Md_shl_out <= (Md_Dout(6 downto 0) & '0');
-------------------------------------------------------------------------------
end structural;
