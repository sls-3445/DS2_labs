------------------------------------------------------------------------------
-- This is the structural description of a neuron for either the hidden or
-- output layers. There is no output activation (rectification) function, but 
-- one like the sigmoid function could be added.
-- (C) April 2019 by Dorin Patru
------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
USE work.sls_package.all;
use work.sls_SSRM_package.all;

------------------------------------------------------------------------------
entity sls_simpleneuron_vhdl is
	port (Reset, Clock, LDmulin, LDmacin, LDz : in std_logic;
			DinA, DinB, biasin : in std_logic_vector(7 downto 0);
			neuronout : out std_logic_vector(7 downto 0));
end sls_simpleneuron_vhdl;
------------------------------------------------------------------------------
architecture structural of sls_simpleneuron_vhdl is
------------------------------------------------------------------------------
-- Internal signals declarations;
------------------------------------------------------------------------------
	signal DmulinA, DmulinB, product_8 : std_logic_vector(7 downto 0);
	signal DaddinA, DaddinB, mac, Dmacout, zin, zout : std_logic_vector(15 downto 0);
	signal product : std_logic_vector(15 downto 0);
	signal cout1, vout1, cout2, vout2 : std_logic;
------------------------------------------------------------------------------
begin
------------------------------------------------------------------------------
-- The two input registers
------------------------------------------------------------------------------
	mulinA : sls_nbit_reg_vhdl generic map (n => 8)
						port map (Reset, Clock, LDmulin, DinA, DmulinA);
	mulinB : sls_nbit_reg_vhdl generic map (n => 8)
						port map (Reset, Clock, LDmulin, DinB, DmulinB);
------------------------------------------------------------------------------
-- This a 16-bit multiplier, i.e. the input operands are each 8-bits wide and 
-- the product 16-bits wide.
-- Replace this with your own multiplier. To match your operand widths, adapt 
-- DmulinA and DmulinB by discarding the most significant bits. To output a 
-- 16-bit product, sign extend your signed product.
------------------------------------------------------------------------------
	mul : sls_16bit_signed_mult_vhdl port map (DmulinA, DmulinB, product);
--	mul : sls_PSRM_vhdl port map (Md_val => DmulinA(3 downto 0), mr_val => DmulinB(3 downto 0), Reset => Reset,
--											Clock => Clock, FP => product_8);
--	product <= (product_8(7) & product_8(7) & product_8(7) & product_8(7) & product_8(7) & 
--				  product_8(7) & product_8(7) & product_8(7) & product_8);
------------------------------------------------------------------------------
-- The MAC accumulator and output register
------------------------------------------------------------------------------
	macinA : sls_nbit_reg_vhdl generic map (n => 16)
						port map (Reset, Clock, LDmacin, product, DaddinA);
	macinB : sls_nbit_reg_vhdl generic map (n => 16)
						port map (Reset, Clock, LDmacin, mac, DaddinB);
------------------------------------------------------------------------------
-- The MAC adder
------------------------------------------------------------------------------
	add1 : sls_16bit_signed_add_vhdl port map (DaddinA, DaddinB, cout1, vout1, mac);
------------------------------------------------------------------------------
-- The MAC accumulator
------------------------------------------------------------------------------
	macinC : sls_nbit_reg_vhdl generic map (n => 16)
						port map (Reset, Clock, LDmacin, mac, Dmacout);
------------------------------------------------------------------------------
-- The BIAS adder
------------------------------------------------------------------------------
--	biasinadjusted <= (biasin(15) & biasin(15) & biasin(15) & biasin(15) & 
--						biasin(15) & biasin(15) & biasin(15) & biasin(15) &
	--						biasin & "00000000"); 
	add2 : sls_16bit_signed_add_vhdl 
						port map (Dmacout, "0000000000000000", cout2, vout2, zin);
------------------------------------------------------------------------------
-- The RAW value output register
------------------------------------------------------------------------------
	zreg : sls_nbit_reg_vhdl generic map (n => 16)
						port map (Reset, Clock, LDz, zin, zout);
------------------------------------------------------------------------------
-- No activation function (rectification/sigmoid) is used.
------------------------------------------------------------------------------
	neuronout <= zout(7 downto 0);
------------------------------------------------------------------------------
end structural;